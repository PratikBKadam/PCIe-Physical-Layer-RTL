module datapath();
endmodule