module LTSSM(input , output );
endmodule
