module tb;
reg clk,rst;
reg [63:0] data_in_LTSSM;
reg [31:0] data_in_DLL;
reg TLP_sent,DLLP_sent,nullified_TLP_sent,framer_en;
wire [7:0] data_1,data_2,data_3,data_4;
wire sender_error_LTSSM,sender_error_DLL;
frame_generator dut(.clk(clk),.rst(rst),.data_in_LTSSM(data_in_LTSSM),.data_1(data_1),.data_2(data_2),.data_3(data_3),.data_4(data_4),
.sender_error_LTSSM(sender_error_LTSSM),.data_in_DLL(data_in_DLL),.TLP_sent(TLP_sent),.DLLP_sent(DLLP_sent),
.nullified_TLP_sent(nullified_TLP_sent),.framer_en(framer_en),.sender_error_DLL(sender_error_DLL));
initial begin
clk=1;
forever #5 clk=~clk;
end
// {TS1_OS,TS2_OS,EIOS,EIEOS,FTS}=buffer[23:19];
// data=buffer[63:24]
// number=buffer[15:0]
initial begin
$monitor("time=%0t, data in LTSSM=0x%0b,\ndata in DLL=0x%0b,\nTLP sent=0x%0b,DLLP sent=0x%0b,nullified TLP sent=0x%0b,framer en=0x%0b,\n data 1=0x%0b,data 2=0x%0b,data 3=0x%0b,data 4=0x%0b ",$time,data_in_LTSSM,data_in_DLL,TLP_sent,DLLP_sent,nullified_TLP_sent,framer_en,data_1,data_2,data_3,data_4);
rst=1'b0;
data_in_LTSSM<=64'h0;
data_in_DLL<=32'h0;
{TLP_sent,DLLP_sent}=2'b0;
framer_en=1'b0;
nullified_TLP_sent=1'b0;
#10;
rst=1'b1;
data_in_LTSSM={8'd1,8'd2,8'd3,8'd4,8'h5,8'b10000000,16'h1};
#10;
data_in_LTSSM=64'h0;
#40;
data_in_LTSSM={8'd1,8'd2,8'd3,8'd4,8'h5,8'b01000000,16'h2};
#10;
data_in_LTSSM=64'h0;
#80;
data_in_LTSSM={8'd1,8'd2,8'd3,8'd4,8'h5,8'b00100000,16'h3};
#10;
data_in_LTSSM=64'h0;
#80;
data_in_LTSSM={8'd1,8'd2,8'd3,8'd4,8'h5,8'b00100001,16'h4};
#10;
data_in_LTSSM=64'h0;
#80;
data_in_LTSSM={8'd1,8'd2,8'd3,8'd4,8'h5,8'b00010000,16'h2};
#10;
data_in_LTSSM=64'h0;
#80;
data_in_LTSSM={8'd1,8'd2,8'd3,8'd4,8'h5,8'b00001000,16'h5};
#10;
data_in_LTSSM=64'h0;
#80;
data_in_LTSSM={8'd1,8'd2,8'd3,8'd4,8'h5,8'b00001001,16'h6};
#10;
data_in_LTSSM=64'h0;
#80;
{TLP_sent,DLLP_sent}=2'b10;
framer_en=1'b0;
data_in_DLL={8'd1,8'd2,8'd3,8'd4};
#10;
rst=1'b1;
{TLP_sent,DLLP_sent}=2'b10;
framer_en=1'b1;
data_in_DLL={8'd5,8'd6,8'd7,8'd8};
#10;
rst=1'b1;
{TLP_sent,DLLP_sent}=2'b10;
framer_en=1'b1;
data_in_DLL={8'd9,8'd10,8'd11,8'd12};
#10;
rst=1'b1;
{TLP_sent,DLLP_sent}=2'b10;
framer_en=1'b1;
data_in_DLL={8'd13,8'd14,8'h0,8'h0};
#10;
{TLP_sent,DLLP_sent}=2'b0;
#10;
framer_en=1'b0;
#10;

{TLP_sent,DLLP_sent}=2'b0;
framer_en=1'b0;
data_in_DLL=32'h0;
#10;
rst=1'b1;
{TLP_sent,DLLP_sent}=2'b01;
framer_en=1'b0;
data_in_DLL={8'd1,8'd2,8'd3,8'd4};
#10;
rst=1'b1;
{TLP_sent,DLLP_sent}=2'b01;
framer_en=1'b1;
data_in_DLL={8'd5,8'd6,8'd7,8'd8};
#10;
rst=1'b1;
{TLP_sent,DLLP_sent}=2'b01;
framer_en=1'b1;
data_in_DLL={8'd9,8'd10,8'h0,8'h0};
#10;
{TLP_sent,DLLP_sent}=2'b0;
#10;
framer_en=1'b0;
#10;

{TLP_sent,DLLP_sent}=2'b00;
framer_en=1'b0;
data_in_DLL=32'h0;
#10;
rst=1'b1;
{TLP_sent,DLLP_sent}=2'b10;
framer_en=1'b0;
data_in_DLL={8'd1,8'd2,8'd3,8'd4};
#10;
rst=1'b1;
{TLP_sent,DLLP_sent}=2'b10;
framer_en=1'b1;
data_in_DLL={8'd5,8'd6,8'd7,8'd8};
#10;
rst=1'b1;
{TLP_sent,DLLP_sent}=2'b10;
framer_en=1'b1;
data_in_DLL={8'd9,8'd10,8'd11,8'd12};
#10;
rst=1'b1;
{TLP_sent,DLLP_sent}=2'b10;
framer_en=1'b1;
data_in_DLL={8'd13,8'd14,8'd0,8'd0};
#10;
{TLP_sent,DLLP_sent}=2'b0;
nullified_TLP_sent=1'b1;
#10;
nullified_TLP_sent=1'b0;
framer_en=1'b0;
#10;
data_in_LTSSM={8'd1,8'd2,8'd3,8'd4,8'h5,8'b10000000,16'h1};
#10;
data_in_LTSSM=64'h0;
#40;
data_in_LTSSM={8'd1,8'd2,8'd3,8'd4,8'h5,8'b01000000,16'h2};
#10;
data_in_LTSSM=64'h0;
#80;
data_in_LTSSM={8'd1,8'd2,8'd3,8'd4,8'h5,8'b00100000,16'h3};
#10;
data_in_LTSSM=64'h0;
#80;
data_in_LTSSM={8'd1,8'd2,8'd3,8'd4,8'h5,8'b00100001,16'h4};
#10;
data_in_LTSSM=64'h0;
#80;
data_in_LTSSM={8'd1,8'd2,8'd3,8'd4,8'h5,8'b00010000,16'h2};
#10;
data_in_LTSSM=64'h0;
#80;
data_in_LTSSM={8'd1,8'd2,8'd3,8'd4,8'h5,8'b00001000,16'h5};
#10;
data_in_LTSSM=64'h0;
#80;
data_in_LTSSM={8'd1,8'd2,8'd3,8'd4,8'h5,8'b00001001,16'h6};
#10;
data_in_LTSSM=64'h0;
#80;
end
endmodule